/******************************************************************************
 ** Logisim-evolution goes FPGA automatic generated Verilog code             **
 ** https://github.com/logisim-evolution/                                    **
 **                                                                          **
 ** Component : srlShift                                                     **
 **                                                                          **
 *****************************************************************************/

module srlShift( in1,
                 out1,
                 shift );

   /*******************************************************************************
   ** The inputs are defined here                                                **
   *******************************************************************************/
   input [31:0] in1;
   input [4:0]  shift;

   /*******************************************************************************
   ** The outputs are defined here                                               **
   *******************************************************************************/
   output [31:0] out1;

   /*******************************************************************************
   ** The wires are defined here                                                 **
   *******************************************************************************/
   wire [31:0] s_logisimBus11;
   wire [31:0] s_logisimBus18;
   wire [31:0] s_logisimBus25;
   wire [31:0] s_logisimBus26;
   wire [31:0] s_logisimBus30;
   wire [31:0] s_logisimBus31;
   wire [31:0] s_logisimBus33;
   wire [31:0] s_logisimBus36;
   wire [31:0] s_logisimBus38;
   wire [31:0] s_logisimBus39;
   wire [31:0] s_logisimBus41;
   wire [31:0] s_logisimBus42;
   wire [31:0] s_logisimBus43;
   wire [31:0] s_logisimBus45;
   wire [31:0] s_logisimBus47;
   wire [31:0] s_logisimBus48;
   wire [31:0] s_logisimBus49;
   wire [31:0] s_logisimBus50;
   wire [31:0] s_logisimBus51;
   wire [31:0] s_logisimBus52;
   wire [31:0] s_logisimBus53;
   wire [31:0] s_logisimBus54;
   wire [31:0] s_logisimBus55;
   wire [31:0] s_logisimBus56;
   wire [31:0] s_logisimBus57;
   wire [31:0] s_logisimBus58;
   wire [31:0] s_logisimBus59;
   wire [31:0] s_logisimBus60;
   wire [31:0] s_logisimBus61;
   wire [31:0] s_logisimBus62;
   wire [31:0] s_logisimBus63;
   wire [31:0] s_logisimBus64;
   wire [31:0] s_logisimBus65;
   wire [4:0]  s_logisimBus9;
   wire        s_logisimNet0;
   wire        s_logisimNet1;
   wire        s_logisimNet10;
   wire        s_logisimNet12;
   wire        s_logisimNet13;
   wire        s_logisimNet14;
   wire        s_logisimNet15;
   wire        s_logisimNet16;
   wire        s_logisimNet17;
   wire        s_logisimNet19;
   wire        s_logisimNet2;
   wire        s_logisimNet20;
   wire        s_logisimNet21;
   wire        s_logisimNet22;
   wire        s_logisimNet23;
   wire        s_logisimNet24;
   wire        s_logisimNet27;
   wire        s_logisimNet28;
   wire        s_logisimNet29;
   wire        s_logisimNet3;
   wire        s_logisimNet32;
   wire        s_logisimNet34;
   wire        s_logisimNet35;
   wire        s_logisimNet37;
   wire        s_logisimNet4;
   wire        s_logisimNet40;
   wire        s_logisimNet44;
   wire        s_logisimNet46;
   wire        s_logisimNet5;
   wire        s_logisimNet6;
   wire        s_logisimNet7;
   wire        s_logisimNet8;

   /*******************************************************************************
   ** The module functionality is described here                                 **
   *******************************************************************************/

   /*******************************************************************************
   ** Here all wiring is defined                                                 **
   *******************************************************************************/
   assign s_logisimBus11[0]  = s_logisimNet46;
   assign s_logisimBus11[10] = s_logisimNet5;
   assign s_logisimBus11[11] = s_logisimNet32;
   assign s_logisimBus11[12] = s_logisimNet13;
   assign s_logisimBus11[13] = s_logisimNet27;
   assign s_logisimBus11[14] = s_logisimNet6;
   assign s_logisimBus11[15] = s_logisimNet3;
   assign s_logisimBus11[16] = s_logisimNet17;
   assign s_logisimBus11[17] = s_logisimNet14;
   assign s_logisimBus11[18] = s_logisimNet24;
   assign s_logisimBus11[19] = s_logisimNet4;
   assign s_logisimBus11[1]  = s_logisimNet37;
   assign s_logisimBus11[20] = s_logisimNet22;
   assign s_logisimBus11[21] = s_logisimNet21;
   assign s_logisimBus11[22] = s_logisimNet20;
   assign s_logisimBus11[23] = s_logisimNet7;
   assign s_logisimBus11[24] = s_logisimNet2;
   assign s_logisimBus11[25] = s_logisimNet23;
   assign s_logisimBus11[26] = s_logisimNet0;
   assign s_logisimBus11[27] = s_logisimNet19;
   assign s_logisimBus11[28] = s_logisimNet16;
   assign s_logisimBus11[29] = s_logisimNet8;
   assign s_logisimBus11[2]  = s_logisimNet35;
   assign s_logisimBus11[30] = s_logisimNet1;
   assign s_logisimBus11[31] = s_logisimNet1;
   assign s_logisimBus11[3]  = s_logisimNet44;
   assign s_logisimBus11[4]  = s_logisimNet29;
   assign s_logisimBus11[5]  = s_logisimNet15;
   assign s_logisimBus11[6]  = s_logisimNet34;
   assign s_logisimBus11[7]  = s_logisimNet12;
   assign s_logisimBus11[8]  = s_logisimNet10;
   assign s_logisimBus11[9]  = s_logisimNet28;
   assign s_logisimBus18[0]  = s_logisimNet32;
   assign s_logisimBus18[10] = s_logisimNet21;
   assign s_logisimBus18[11] = s_logisimNet20;
   assign s_logisimBus18[12] = s_logisimNet7;
   assign s_logisimBus18[13] = s_logisimNet2;
   assign s_logisimBus18[14] = s_logisimNet23;
   assign s_logisimBus18[15] = s_logisimNet0;
   assign s_logisimBus18[16] = s_logisimNet19;
   assign s_logisimBus18[17] = s_logisimNet16;
   assign s_logisimBus18[18] = s_logisimNet8;
   assign s_logisimBus18[19] = s_logisimNet1;
   assign s_logisimBus18[1]  = s_logisimNet13;
   assign s_logisimBus18[20] = s_logisimNet1;
   assign s_logisimBus18[21] = s_logisimNet1;
   assign s_logisimBus18[22] = s_logisimNet1;
   assign s_logisimBus18[23] = s_logisimNet1;
   assign s_logisimBus18[24] = s_logisimNet1;
   assign s_logisimBus18[25] = s_logisimNet1;
   assign s_logisimBus18[26] = s_logisimNet1;
   assign s_logisimBus18[27] = s_logisimNet1;
   assign s_logisimBus18[28] = s_logisimNet1;
   assign s_logisimBus18[29] = s_logisimNet1;
   assign s_logisimBus18[2]  = s_logisimNet27;
   assign s_logisimBus18[30] = s_logisimNet1;
   assign s_logisimBus18[31] = s_logisimNet1;
   assign s_logisimBus18[3]  = s_logisimNet6;
   assign s_logisimBus18[4]  = s_logisimNet3;
   assign s_logisimBus18[5]  = s_logisimNet17;
   assign s_logisimBus18[6]  = s_logisimNet14;
   assign s_logisimBus18[7]  = s_logisimNet24;
   assign s_logisimBus18[8]  = s_logisimNet4;
   assign s_logisimBus18[9]  = s_logisimNet22;
   assign s_logisimBus26[0]  = s_logisimNet37;
   assign s_logisimBus26[10] = s_logisimNet32;
   assign s_logisimBus26[11] = s_logisimNet13;
   assign s_logisimBus26[12] = s_logisimNet27;
   assign s_logisimBus26[13] = s_logisimNet6;
   assign s_logisimBus26[14] = s_logisimNet3;
   assign s_logisimBus26[15] = s_logisimNet17;
   assign s_logisimBus26[16] = s_logisimNet14;
   assign s_logisimBus26[17] = s_logisimNet24;
   assign s_logisimBus26[18] = s_logisimNet4;
   assign s_logisimBus26[19] = s_logisimNet22;
   assign s_logisimBus26[1]  = s_logisimNet35;
   assign s_logisimBus26[20] = s_logisimNet21;
   assign s_logisimBus26[21] = s_logisimNet20;
   assign s_logisimBus26[22] = s_logisimNet7;
   assign s_logisimBus26[23] = s_logisimNet2;
   assign s_logisimBus26[24] = s_logisimNet23;
   assign s_logisimBus26[25] = s_logisimNet0;
   assign s_logisimBus26[26] = s_logisimNet19;
   assign s_logisimBus26[27] = s_logisimNet16;
   assign s_logisimBus26[28] = s_logisimNet8;
   assign s_logisimBus26[29] = s_logisimNet1;
   assign s_logisimBus26[2]  = s_logisimNet44;
   assign s_logisimBus26[30] = s_logisimNet1;
   assign s_logisimBus26[31] = s_logisimNet1;
   assign s_logisimBus26[3]  = s_logisimNet29;
   assign s_logisimBus26[4]  = s_logisimNet15;
   assign s_logisimBus26[5]  = s_logisimNet34;
   assign s_logisimBus26[6]  = s_logisimNet12;
   assign s_logisimBus26[7]  = s_logisimNet10;
   assign s_logisimBus26[8]  = s_logisimNet28;
   assign s_logisimBus26[9]  = s_logisimNet5;
   assign s_logisimBus30[0]  = s_logisimNet0;
   assign s_logisimBus30[10] = s_logisimNet1;
   assign s_logisimBus30[11] = s_logisimNet1;
   assign s_logisimBus30[12] = s_logisimNet1;
   assign s_logisimBus30[13] = s_logisimNet1;
   assign s_logisimBus30[14] = s_logisimNet1;
   assign s_logisimBus30[15] = s_logisimNet1;
   assign s_logisimBus30[16] = s_logisimNet1;
   assign s_logisimBus30[17] = s_logisimNet1;
   assign s_logisimBus30[18] = s_logisimNet1;
   assign s_logisimBus30[19] = s_logisimNet1;
   assign s_logisimBus30[1]  = s_logisimNet19;
   assign s_logisimBus30[20] = s_logisimNet1;
   assign s_logisimBus30[21] = s_logisimNet1;
   assign s_logisimBus30[22] = s_logisimNet1;
   assign s_logisimBus30[23] = s_logisimNet1;
   assign s_logisimBus30[24] = s_logisimNet1;
   assign s_logisimBus30[25] = s_logisimNet1;
   assign s_logisimBus30[26] = s_logisimNet1;
   assign s_logisimBus30[27] = s_logisimNet1;
   assign s_logisimBus30[28] = s_logisimNet1;
   assign s_logisimBus30[29] = s_logisimNet1;
   assign s_logisimBus30[2]  = s_logisimNet16;
   assign s_logisimBus30[30] = s_logisimNet1;
   assign s_logisimBus30[31] = s_logisimNet1;
   assign s_logisimBus30[3]  = s_logisimNet8;
   assign s_logisimBus30[4]  = s_logisimNet1;
   assign s_logisimBus30[5]  = s_logisimNet1;
   assign s_logisimBus30[6]  = s_logisimNet1;
   assign s_logisimBus30[7]  = s_logisimNet1;
   assign s_logisimBus30[8]  = s_logisimNet1;
   assign s_logisimBus30[9]  = s_logisimNet1;
   assign s_logisimBus31[0]  = s_logisimNet19;
   assign s_logisimBus31[10] = s_logisimNet1;
   assign s_logisimBus31[11] = s_logisimNet1;
   assign s_logisimBus31[12] = s_logisimNet1;
   assign s_logisimBus31[13] = s_logisimNet1;
   assign s_logisimBus31[14] = s_logisimNet1;
   assign s_logisimBus31[15] = s_logisimNet1;
   assign s_logisimBus31[16] = s_logisimNet1;
   assign s_logisimBus31[17] = s_logisimNet1;
   assign s_logisimBus31[18] = s_logisimNet1;
   assign s_logisimBus31[19] = s_logisimNet1;
   assign s_logisimBus31[1]  = s_logisimNet16;
   assign s_logisimBus31[20] = s_logisimNet1;
   assign s_logisimBus31[21] = s_logisimNet1;
   assign s_logisimBus31[22] = s_logisimNet1;
   assign s_logisimBus31[23] = s_logisimNet1;
   assign s_logisimBus31[24] = s_logisimNet1;
   assign s_logisimBus31[25] = s_logisimNet1;
   assign s_logisimBus31[26] = s_logisimNet1;
   assign s_logisimBus31[27] = s_logisimNet1;
   assign s_logisimBus31[28] = s_logisimNet1;
   assign s_logisimBus31[29] = s_logisimNet1;
   assign s_logisimBus31[2]  = s_logisimNet8;
   assign s_logisimBus31[30] = s_logisimNet1;
   assign s_logisimBus31[31] = s_logisimNet1;
   assign s_logisimBus31[3]  = s_logisimNet1;
   assign s_logisimBus31[4]  = s_logisimNet1;
   assign s_logisimBus31[5]  = s_logisimNet1;
   assign s_logisimBus31[6]  = s_logisimNet1;
   assign s_logisimBus31[7]  = s_logisimNet1;
   assign s_logisimBus31[8]  = s_logisimNet1;
   assign s_logisimBus31[9]  = s_logisimNet1;
   assign s_logisimBus33[0]  = s_logisimNet5;
   assign s_logisimBus33[10] = s_logisimNet22;
   assign s_logisimBus33[11] = s_logisimNet21;
   assign s_logisimBus33[12] = s_logisimNet20;
   assign s_logisimBus33[13] = s_logisimNet7;
   assign s_logisimBus33[14] = s_logisimNet2;
   assign s_logisimBus33[15] = s_logisimNet23;
   assign s_logisimBus33[16] = s_logisimNet0;
   assign s_logisimBus33[17] = s_logisimNet19;
   assign s_logisimBus33[18] = s_logisimNet16;
   assign s_logisimBus33[19] = s_logisimNet8;
   assign s_logisimBus33[1]  = s_logisimNet32;
   assign s_logisimBus33[20] = s_logisimNet1;
   assign s_logisimBus33[21] = s_logisimNet1;
   assign s_logisimBus33[22] = s_logisimNet1;
   assign s_logisimBus33[23] = s_logisimNet1;
   assign s_logisimBus33[24] = s_logisimNet1;
   assign s_logisimBus33[25] = s_logisimNet1;
   assign s_logisimBus33[26] = s_logisimNet1;
   assign s_logisimBus33[27] = s_logisimNet1;
   assign s_logisimBus33[28] = s_logisimNet1;
   assign s_logisimBus33[29] = s_logisimNet1;
   assign s_logisimBus33[2]  = s_logisimNet13;
   assign s_logisimBus33[30] = s_logisimNet1;
   assign s_logisimBus33[31] = s_logisimNet1;
   assign s_logisimBus33[3]  = s_logisimNet27;
   assign s_logisimBus33[4]  = s_logisimNet6;
   assign s_logisimBus33[5]  = s_logisimNet3;
   assign s_logisimBus33[6]  = s_logisimNet17;
   assign s_logisimBus33[7]  = s_logisimNet14;
   assign s_logisimBus33[8]  = s_logisimNet24;
   assign s_logisimBus33[9]  = s_logisimNet4;
   assign s_logisimBus36[0]  = s_logisimNet24;
   assign s_logisimBus36[10] = s_logisimNet16;
   assign s_logisimBus36[11] = s_logisimNet8;
   assign s_logisimBus36[12] = s_logisimNet1;
   assign s_logisimBus36[13] = s_logisimNet1;
   assign s_logisimBus36[14] = s_logisimNet1;
   assign s_logisimBus36[15] = s_logisimNet1;
   assign s_logisimBus36[16] = s_logisimNet1;
   assign s_logisimBus36[17] = s_logisimNet1;
   assign s_logisimBus36[18] = s_logisimNet1;
   assign s_logisimBus36[19] = s_logisimNet1;
   assign s_logisimBus36[1]  = s_logisimNet4;
   assign s_logisimBus36[20] = s_logisimNet1;
   assign s_logisimBus36[21] = s_logisimNet1;
   assign s_logisimBus36[22] = s_logisimNet1;
   assign s_logisimBus36[23] = s_logisimNet1;
   assign s_logisimBus36[24] = s_logisimNet1;
   assign s_logisimBus36[25] = s_logisimNet1;
   assign s_logisimBus36[26] = s_logisimNet1;
   assign s_logisimBus36[27] = s_logisimNet1;
   assign s_logisimBus36[28] = s_logisimNet1;
   assign s_logisimBus36[29] = s_logisimNet1;
   assign s_logisimBus36[2]  = s_logisimNet22;
   assign s_logisimBus36[30] = s_logisimNet1;
   assign s_logisimBus36[31] = s_logisimNet1;
   assign s_logisimBus36[3]  = s_logisimNet21;
   assign s_logisimBus36[4]  = s_logisimNet20;
   assign s_logisimBus36[5]  = s_logisimNet7;
   assign s_logisimBus36[6]  = s_logisimNet2;
   assign s_logisimBus36[7]  = s_logisimNet23;
   assign s_logisimBus36[8]  = s_logisimNet0;
   assign s_logisimBus36[9]  = s_logisimNet19;
   assign s_logisimBus38[0]  = s_logisimNet16;
   assign s_logisimBus38[10] = s_logisimNet1;
   assign s_logisimBus38[11] = s_logisimNet1;
   assign s_logisimBus38[12] = s_logisimNet1;
   assign s_logisimBus38[13] = s_logisimNet1;
   assign s_logisimBus38[14] = s_logisimNet1;
   assign s_logisimBus38[15] = s_logisimNet1;
   assign s_logisimBus38[16] = s_logisimNet1;
   assign s_logisimBus38[17] = s_logisimNet1;
   assign s_logisimBus38[18] = s_logisimNet1;
   assign s_logisimBus38[19] = s_logisimNet1;
   assign s_logisimBus38[1]  = s_logisimNet8;
   assign s_logisimBus38[20] = s_logisimNet1;
   assign s_logisimBus38[21] = s_logisimNet1;
   assign s_logisimBus38[22] = s_logisimNet1;
   assign s_logisimBus38[23] = s_logisimNet1;
   assign s_logisimBus38[24] = s_logisimNet1;
   assign s_logisimBus38[25] = s_logisimNet1;
   assign s_logisimBus38[26] = s_logisimNet1;
   assign s_logisimBus38[27] = s_logisimNet1;
   assign s_logisimBus38[28] = s_logisimNet1;
   assign s_logisimBus38[29] = s_logisimNet1;
   assign s_logisimBus38[2]  = s_logisimNet1;
   assign s_logisimBus38[30] = s_logisimNet1;
   assign s_logisimBus38[31] = s_logisimNet1;
   assign s_logisimBus38[3]  = s_logisimNet1;
   assign s_logisimBus38[4]  = s_logisimNet1;
   assign s_logisimBus38[5]  = s_logisimNet1;
   assign s_logisimBus38[6]  = s_logisimNet1;
   assign s_logisimBus38[7]  = s_logisimNet1;
   assign s_logisimBus38[8]  = s_logisimNet1;
   assign s_logisimBus38[9]  = s_logisimNet1;
   assign s_logisimBus39[0]  = s_logisimNet28;
   assign s_logisimBus39[10] = s_logisimNet4;
   assign s_logisimBus39[11] = s_logisimNet22;
   assign s_logisimBus39[12] = s_logisimNet21;
   assign s_logisimBus39[13] = s_logisimNet20;
   assign s_logisimBus39[14] = s_logisimNet7;
   assign s_logisimBus39[15] = s_logisimNet2;
   assign s_logisimBus39[16] = s_logisimNet23;
   assign s_logisimBus39[17] = s_logisimNet0;
   assign s_logisimBus39[18] = s_logisimNet19;
   assign s_logisimBus39[19] = s_logisimNet16;
   assign s_logisimBus39[1]  = s_logisimNet5;
   assign s_logisimBus39[20] = s_logisimNet8;
   assign s_logisimBus39[21] = s_logisimNet1;
   assign s_logisimBus39[22] = s_logisimNet1;
   assign s_logisimBus39[23] = s_logisimNet1;
   assign s_logisimBus39[24] = s_logisimNet1;
   assign s_logisimBus39[25] = s_logisimNet1;
   assign s_logisimBus39[26] = s_logisimNet1;
   assign s_logisimBus39[27] = s_logisimNet1;
   assign s_logisimBus39[28] = s_logisimNet1;
   assign s_logisimBus39[29] = s_logisimNet1;
   assign s_logisimBus39[2]  = s_logisimNet32;
   assign s_logisimBus39[30] = s_logisimNet1;
   assign s_logisimBus39[31] = s_logisimNet1;
   assign s_logisimBus39[3]  = s_logisimNet13;
   assign s_logisimBus39[4]  = s_logisimNet27;
   assign s_logisimBus39[5]  = s_logisimNet6;
   assign s_logisimBus39[6]  = s_logisimNet3;
   assign s_logisimBus39[7]  = s_logisimNet17;
   assign s_logisimBus39[8]  = s_logisimNet14;
   assign s_logisimBus39[9]  = s_logisimNet24;
   assign s_logisimBus41[0]  = s_logisimNet15;
   assign s_logisimBus41[10] = s_logisimNet3;
   assign s_logisimBus41[11] = s_logisimNet17;
   assign s_logisimBus41[12] = s_logisimNet14;
   assign s_logisimBus41[13] = s_logisimNet24;
   assign s_logisimBus41[14] = s_logisimNet4;
   assign s_logisimBus41[15] = s_logisimNet22;
   assign s_logisimBus41[16] = s_logisimNet21;
   assign s_logisimBus41[17] = s_logisimNet20;
   assign s_logisimBus41[18] = s_logisimNet7;
   assign s_logisimBus41[19] = s_logisimNet2;
   assign s_logisimBus41[1]  = s_logisimNet34;
   assign s_logisimBus41[20] = s_logisimNet23;
   assign s_logisimBus41[21] = s_logisimNet0;
   assign s_logisimBus41[22] = s_logisimNet19;
   assign s_logisimBus41[23] = s_logisimNet16;
   assign s_logisimBus41[24] = s_logisimNet8;
   assign s_logisimBus41[25] = s_logisimNet1;
   assign s_logisimBus41[26] = s_logisimNet1;
   assign s_logisimBus41[27] = s_logisimNet1;
   assign s_logisimBus41[28] = s_logisimNet1;
   assign s_logisimBus41[29] = s_logisimNet1;
   assign s_logisimBus41[2]  = s_logisimNet12;
   assign s_logisimBus41[30] = s_logisimNet1;
   assign s_logisimBus41[31] = s_logisimNet1;
   assign s_logisimBus41[3]  = s_logisimNet10;
   assign s_logisimBus41[4]  = s_logisimNet28;
   assign s_logisimBus41[5]  = s_logisimNet5;
   assign s_logisimBus41[6]  = s_logisimNet32;
   assign s_logisimBus41[7]  = s_logisimNet13;
   assign s_logisimBus41[8]  = s_logisimNet27;
   assign s_logisimBus41[9]  = s_logisimNet6;
   assign s_logisimBus42[0]  = s_logisimNet14;
   assign s_logisimBus42[10] = s_logisimNet19;
   assign s_logisimBus42[11] = s_logisimNet16;
   assign s_logisimBus42[12] = s_logisimNet8;
   assign s_logisimBus42[13] = s_logisimNet1;
   assign s_logisimBus42[14] = s_logisimNet1;
   assign s_logisimBus42[15] = s_logisimNet1;
   assign s_logisimBus42[16] = s_logisimNet1;
   assign s_logisimBus42[17] = s_logisimNet1;
   assign s_logisimBus42[18] = s_logisimNet1;
   assign s_logisimBus42[19] = s_logisimNet1;
   assign s_logisimBus42[1]  = s_logisimNet24;
   assign s_logisimBus42[20] = s_logisimNet1;
   assign s_logisimBus42[21] = s_logisimNet1;
   assign s_logisimBus42[22] = s_logisimNet1;
   assign s_logisimBus42[23] = s_logisimNet1;
   assign s_logisimBus42[24] = s_logisimNet1;
   assign s_logisimBus42[25] = s_logisimNet1;
   assign s_logisimBus42[26] = s_logisimNet1;
   assign s_logisimBus42[27] = s_logisimNet1;
   assign s_logisimBus42[28] = s_logisimNet1;
   assign s_logisimBus42[29] = s_logisimNet1;
   assign s_logisimBus42[2]  = s_logisimNet4;
   assign s_logisimBus42[30] = s_logisimNet1;
   assign s_logisimBus42[31] = s_logisimNet1;
   assign s_logisimBus42[3]  = s_logisimNet22;
   assign s_logisimBus42[4]  = s_logisimNet21;
   assign s_logisimBus42[5]  = s_logisimNet20;
   assign s_logisimBus42[6]  = s_logisimNet7;
   assign s_logisimBus42[7]  = s_logisimNet2;
   assign s_logisimBus42[8]  = s_logisimNet23;
   assign s_logisimBus42[9]  = s_logisimNet0;
   assign s_logisimBus43[0]  = s_logisimNet2;
   assign s_logisimBus43[10] = s_logisimNet1;
   assign s_logisimBus43[11] = s_logisimNet1;
   assign s_logisimBus43[12] = s_logisimNet1;
   assign s_logisimBus43[13] = s_logisimNet1;
   assign s_logisimBus43[14] = s_logisimNet1;
   assign s_logisimBus43[15] = s_logisimNet1;
   assign s_logisimBus43[16] = s_logisimNet1;
   assign s_logisimBus43[17] = s_logisimNet1;
   assign s_logisimBus43[18] = s_logisimNet1;
   assign s_logisimBus43[19] = s_logisimNet1;
   assign s_logisimBus43[1]  = s_logisimNet23;
   assign s_logisimBus43[20] = s_logisimNet1;
   assign s_logisimBus43[21] = s_logisimNet1;
   assign s_logisimBus43[22] = s_logisimNet1;
   assign s_logisimBus43[23] = s_logisimNet1;
   assign s_logisimBus43[24] = s_logisimNet1;
   assign s_logisimBus43[25] = s_logisimNet1;
   assign s_logisimBus43[26] = s_logisimNet1;
   assign s_logisimBus43[27] = s_logisimNet1;
   assign s_logisimBus43[28] = s_logisimNet1;
   assign s_logisimBus43[29] = s_logisimNet1;
   assign s_logisimBus43[2]  = s_logisimNet0;
   assign s_logisimBus43[30] = s_logisimNet1;
   assign s_logisimBus43[31] = s_logisimNet1;
   assign s_logisimBus43[3]  = s_logisimNet19;
   assign s_logisimBus43[4]  = s_logisimNet16;
   assign s_logisimBus43[5]  = s_logisimNet8;
   assign s_logisimBus43[6]  = s_logisimNet1;
   assign s_logisimBus43[7]  = s_logisimNet1;
   assign s_logisimBus43[8]  = s_logisimNet1;
   assign s_logisimBus43[9]  = s_logisimNet1;
   assign s_logisimBus45[0]  = s_logisimNet29;
   assign s_logisimBus45[10] = s_logisimNet6;
   assign s_logisimBus45[11] = s_logisimNet3;
   assign s_logisimBus45[12] = s_logisimNet17;
   assign s_logisimBus45[13] = s_logisimNet14;
   assign s_logisimBus45[14] = s_logisimNet24;
   assign s_logisimBus45[15] = s_logisimNet4;
   assign s_logisimBus45[16] = s_logisimNet22;
   assign s_logisimBus45[17] = s_logisimNet21;
   assign s_logisimBus45[18] = s_logisimNet20;
   assign s_logisimBus45[19] = s_logisimNet7;
   assign s_logisimBus45[1]  = s_logisimNet15;
   assign s_logisimBus45[20] = s_logisimNet2;
   assign s_logisimBus45[21] = s_logisimNet23;
   assign s_logisimBus45[22] = s_logisimNet0;
   assign s_logisimBus45[23] = s_logisimNet19;
   assign s_logisimBus45[24] = s_logisimNet16;
   assign s_logisimBus45[25] = s_logisimNet8;
   assign s_logisimBus45[26] = s_logisimNet1;
   assign s_logisimBus45[27] = s_logisimNet1;
   assign s_logisimBus45[28] = s_logisimNet1;
   assign s_logisimBus45[29] = s_logisimNet1;
   assign s_logisimBus45[2]  = s_logisimNet34;
   assign s_logisimBus45[30] = s_logisimNet1;
   assign s_logisimBus45[31] = s_logisimNet1;
   assign s_logisimBus45[3]  = s_logisimNet12;
   assign s_logisimBus45[4]  = s_logisimNet10;
   assign s_logisimBus45[5]  = s_logisimNet28;
   assign s_logisimBus45[6]  = s_logisimNet5;
   assign s_logisimBus45[7]  = s_logisimNet32;
   assign s_logisimBus45[8]  = s_logisimNet13;
   assign s_logisimBus45[9]  = s_logisimNet27;
   assign s_logisimBus47[0]  = s_logisimNet13;
   assign s_logisimBus47[10] = s_logisimNet20;
   assign s_logisimBus47[11] = s_logisimNet7;
   assign s_logisimBus47[12] = s_logisimNet2;
   assign s_logisimBus47[13] = s_logisimNet23;
   assign s_logisimBus47[14] = s_logisimNet0;
   assign s_logisimBus47[15] = s_logisimNet19;
   assign s_logisimBus47[16] = s_logisimNet16;
   assign s_logisimBus47[17] = s_logisimNet8;
   assign s_logisimBus47[18] = s_logisimNet1;
   assign s_logisimBus47[19] = s_logisimNet1;
   assign s_logisimBus47[1]  = s_logisimNet27;
   assign s_logisimBus47[20] = s_logisimNet1;
   assign s_logisimBus47[21] = s_logisimNet1;
   assign s_logisimBus47[22] = s_logisimNet1;
   assign s_logisimBus47[23] = s_logisimNet1;
   assign s_logisimBus47[24] = s_logisimNet1;
   assign s_logisimBus47[25] = s_logisimNet1;
   assign s_logisimBus47[26] = s_logisimNet1;
   assign s_logisimBus47[27] = s_logisimNet1;
   assign s_logisimBus47[28] = s_logisimNet1;
   assign s_logisimBus47[29] = s_logisimNet1;
   assign s_logisimBus47[2]  = s_logisimNet6;
   assign s_logisimBus47[30] = s_logisimNet1;
   assign s_logisimBus47[31] = s_logisimNet1;
   assign s_logisimBus47[3]  = s_logisimNet3;
   assign s_logisimBus47[4]  = s_logisimNet17;
   assign s_logisimBus47[5]  = s_logisimNet14;
   assign s_logisimBus47[6]  = s_logisimNet24;
   assign s_logisimBus47[7]  = s_logisimNet4;
   assign s_logisimBus47[8]  = s_logisimNet22;
   assign s_logisimBus47[9]  = s_logisimNet21;
   assign s_logisimBus48[0]  = s_logisimNet8;
   assign s_logisimBus48[10] = s_logisimNet1;
   assign s_logisimBus48[11] = s_logisimNet1;
   assign s_logisimBus48[12] = s_logisimNet1;
   assign s_logisimBus48[13] = s_logisimNet1;
   assign s_logisimBus48[14] = s_logisimNet1;
   assign s_logisimBus48[15] = s_logisimNet1;
   assign s_logisimBus48[16] = s_logisimNet1;
   assign s_logisimBus48[17] = s_logisimNet1;
   assign s_logisimBus48[18] = s_logisimNet1;
   assign s_logisimBus48[19] = s_logisimNet1;
   assign s_logisimBus48[1]  = s_logisimNet1;
   assign s_logisimBus48[20] = s_logisimNet1;
   assign s_logisimBus48[21] = s_logisimNet1;
   assign s_logisimBus48[22] = s_logisimNet1;
   assign s_logisimBus48[23] = s_logisimNet1;
   assign s_logisimBus48[24] = s_logisimNet1;
   assign s_logisimBus48[25] = s_logisimNet1;
   assign s_logisimBus48[26] = s_logisimNet1;
   assign s_logisimBus48[27] = s_logisimNet1;
   assign s_logisimBus48[28] = s_logisimNet1;
   assign s_logisimBus48[29] = s_logisimNet1;
   assign s_logisimBus48[2]  = s_logisimNet1;
   assign s_logisimBus48[30] = s_logisimNet1;
   assign s_logisimBus48[31] = s_logisimNet1;
   assign s_logisimBus48[3]  = s_logisimNet1;
   assign s_logisimBus48[4]  = s_logisimNet1;
   assign s_logisimBus48[5]  = s_logisimNet1;
   assign s_logisimBus48[6]  = s_logisimNet1;
   assign s_logisimBus48[7]  = s_logisimNet1;
   assign s_logisimBus48[8]  = s_logisimNet1;
   assign s_logisimBus48[9]  = s_logisimNet1;
   assign s_logisimBus49[0]  = s_logisimNet23;
   assign s_logisimBus49[10] = s_logisimNet1;
   assign s_logisimBus49[11] = s_logisimNet1;
   assign s_logisimBus49[12] = s_logisimNet1;
   assign s_logisimBus49[13] = s_logisimNet1;
   assign s_logisimBus49[14] = s_logisimNet1;
   assign s_logisimBus49[15] = s_logisimNet1;
   assign s_logisimBus49[16] = s_logisimNet1;
   assign s_logisimBus49[17] = s_logisimNet1;
   assign s_logisimBus49[18] = s_logisimNet1;
   assign s_logisimBus49[19] = s_logisimNet1;
   assign s_logisimBus49[1]  = s_logisimNet0;
   assign s_logisimBus49[20] = s_logisimNet1;
   assign s_logisimBus49[21] = s_logisimNet1;
   assign s_logisimBus49[22] = s_logisimNet1;
   assign s_logisimBus49[23] = s_logisimNet1;
   assign s_logisimBus49[24] = s_logisimNet1;
   assign s_logisimBus49[25] = s_logisimNet1;
   assign s_logisimBus49[26] = s_logisimNet1;
   assign s_logisimBus49[27] = s_logisimNet1;
   assign s_logisimBus49[28] = s_logisimNet1;
   assign s_logisimBus49[29] = s_logisimNet1;
   assign s_logisimBus49[2]  = s_logisimNet19;
   assign s_logisimBus49[30] = s_logisimNet1;
   assign s_logisimBus49[31] = s_logisimNet1;
   assign s_logisimBus49[3]  = s_logisimNet16;
   assign s_logisimBus49[4]  = s_logisimNet8;
   assign s_logisimBus49[5]  = s_logisimNet1;
   assign s_logisimBus49[6]  = s_logisimNet1;
   assign s_logisimBus49[7]  = s_logisimNet1;
   assign s_logisimBus49[8]  = s_logisimNet1;
   assign s_logisimBus49[9]  = s_logisimNet1;
   assign s_logisimBus50[0]  = s_logisimNet21;
   assign s_logisimBus50[10] = s_logisimNet1;
   assign s_logisimBus50[11] = s_logisimNet1;
   assign s_logisimBus50[12] = s_logisimNet1;
   assign s_logisimBus50[13] = s_logisimNet1;
   assign s_logisimBus50[14] = s_logisimNet1;
   assign s_logisimBus50[15] = s_logisimNet1;
   assign s_logisimBus50[16] = s_logisimNet1;
   assign s_logisimBus50[17] = s_logisimNet1;
   assign s_logisimBus50[18] = s_logisimNet1;
   assign s_logisimBus50[19] = s_logisimNet1;
   assign s_logisimBus50[1]  = s_logisimNet20;
   assign s_logisimBus50[20] = s_logisimNet1;
   assign s_logisimBus50[21] = s_logisimNet1;
   assign s_logisimBus50[22] = s_logisimNet1;
   assign s_logisimBus50[23] = s_logisimNet1;
   assign s_logisimBus50[24] = s_logisimNet1;
   assign s_logisimBus50[25] = s_logisimNet1;
   assign s_logisimBus50[26] = s_logisimNet1;
   assign s_logisimBus50[27] = s_logisimNet1;
   assign s_logisimBus50[28] = s_logisimNet1;
   assign s_logisimBus50[29] = s_logisimNet1;
   assign s_logisimBus50[2]  = s_logisimNet7;
   assign s_logisimBus50[30] = s_logisimNet1;
   assign s_logisimBus50[31] = s_logisimNet1;
   assign s_logisimBus50[3]  = s_logisimNet2;
   assign s_logisimBus50[4]  = s_logisimNet23;
   assign s_logisimBus50[5]  = s_logisimNet0;
   assign s_logisimBus50[6]  = s_logisimNet19;
   assign s_logisimBus50[7]  = s_logisimNet16;
   assign s_logisimBus50[8]  = s_logisimNet8;
   assign s_logisimBus50[9]  = s_logisimNet1;
   assign s_logisimBus51[0]  = s_logisimNet34;
   assign s_logisimBus51[10] = s_logisimNet17;
   assign s_logisimBus51[11] = s_logisimNet14;
   assign s_logisimBus51[12] = s_logisimNet24;
   assign s_logisimBus51[13] = s_logisimNet4;
   assign s_logisimBus51[14] = s_logisimNet22;
   assign s_logisimBus51[15] = s_logisimNet21;
   assign s_logisimBus51[16] = s_logisimNet20;
   assign s_logisimBus51[17] = s_logisimNet7;
   assign s_logisimBus51[18] = s_logisimNet2;
   assign s_logisimBus51[19] = s_logisimNet23;
   assign s_logisimBus51[1]  = s_logisimNet12;
   assign s_logisimBus51[20] = s_logisimNet0;
   assign s_logisimBus51[21] = s_logisimNet19;
   assign s_logisimBus51[22] = s_logisimNet16;
   assign s_logisimBus51[23] = s_logisimNet8;
   assign s_logisimBus51[24] = s_logisimNet1;
   assign s_logisimBus51[25] = s_logisimNet1;
   assign s_logisimBus51[26] = s_logisimNet1;
   assign s_logisimBus51[27] = s_logisimNet1;
   assign s_logisimBus51[28] = s_logisimNet1;
   assign s_logisimBus51[29] = s_logisimNet1;
   assign s_logisimBus51[2]  = s_logisimNet10;
   assign s_logisimBus51[30] = s_logisimNet1;
   assign s_logisimBus51[31] = s_logisimNet1;
   assign s_logisimBus51[3]  = s_logisimNet28;
   assign s_logisimBus51[4]  = s_logisimNet5;
   assign s_logisimBus51[5]  = s_logisimNet32;
   assign s_logisimBus51[6]  = s_logisimNet13;
   assign s_logisimBus51[7]  = s_logisimNet27;
   assign s_logisimBus51[8]  = s_logisimNet6;
   assign s_logisimBus51[9]  = s_logisimNet3;
   assign s_logisimBus52[0]  = s_logisimNet6;
   assign s_logisimBus52[10] = s_logisimNet2;
   assign s_logisimBus52[11] = s_logisimNet23;
   assign s_logisimBus52[12] = s_logisimNet0;
   assign s_logisimBus52[13] = s_logisimNet19;
   assign s_logisimBus52[14] = s_logisimNet16;
   assign s_logisimBus52[15] = s_logisimNet8;
   assign s_logisimBus52[16] = s_logisimNet1;
   assign s_logisimBus52[17] = s_logisimNet1;
   assign s_logisimBus52[18] = s_logisimNet1;
   assign s_logisimBus52[19] = s_logisimNet1;
   assign s_logisimBus52[1]  = s_logisimNet3;
   assign s_logisimBus52[20] = s_logisimNet1;
   assign s_logisimBus52[21] = s_logisimNet1;
   assign s_logisimBus52[22] = s_logisimNet1;
   assign s_logisimBus52[23] = s_logisimNet1;
   assign s_logisimBus52[24] = s_logisimNet1;
   assign s_logisimBus52[25] = s_logisimNet1;
   assign s_logisimBus52[26] = s_logisimNet1;
   assign s_logisimBus52[27] = s_logisimNet1;
   assign s_logisimBus52[28] = s_logisimNet1;
   assign s_logisimBus52[29] = s_logisimNet1;
   assign s_logisimBus52[2]  = s_logisimNet17;
   assign s_logisimBus52[30] = s_logisimNet1;
   assign s_logisimBus52[31] = s_logisimNet1;
   assign s_logisimBus52[3]  = s_logisimNet14;
   assign s_logisimBus52[4]  = s_logisimNet24;
   assign s_logisimBus52[5]  = s_logisimNet4;
   assign s_logisimBus52[6]  = s_logisimNet22;
   assign s_logisimBus52[7]  = s_logisimNet21;
   assign s_logisimBus52[8]  = s_logisimNet20;
   assign s_logisimBus52[9]  = s_logisimNet7;
   assign s_logisimBus53[0]  = s_logisimNet10;
   assign s_logisimBus53[10] = s_logisimNet24;
   assign s_logisimBus53[11] = s_logisimNet4;
   assign s_logisimBus53[12] = s_logisimNet22;
   assign s_logisimBus53[13] = s_logisimNet21;
   assign s_logisimBus53[14] = s_logisimNet20;
   assign s_logisimBus53[15] = s_logisimNet7;
   assign s_logisimBus53[16] = s_logisimNet2;
   assign s_logisimBus53[17] = s_logisimNet23;
   assign s_logisimBus53[18] = s_logisimNet0;
   assign s_logisimBus53[19] = s_logisimNet19;
   assign s_logisimBus53[1]  = s_logisimNet28;
   assign s_logisimBus53[20] = s_logisimNet16;
   assign s_logisimBus53[21] = s_logisimNet8;
   assign s_logisimBus53[22] = s_logisimNet1;
   assign s_logisimBus53[23] = s_logisimNet1;
   assign s_logisimBus53[24] = s_logisimNet1;
   assign s_logisimBus53[25] = s_logisimNet1;
   assign s_logisimBus53[26] = s_logisimNet1;
   assign s_logisimBus53[27] = s_logisimNet1;
   assign s_logisimBus53[28] = s_logisimNet1;
   assign s_logisimBus53[29] = s_logisimNet1;
   assign s_logisimBus53[2]  = s_logisimNet5;
   assign s_logisimBus53[30] = s_logisimNet1;
   assign s_logisimBus53[31] = s_logisimNet1;
   assign s_logisimBus53[3]  = s_logisimNet32;
   assign s_logisimBus53[4]  = s_logisimNet13;
   assign s_logisimBus53[5]  = s_logisimNet27;
   assign s_logisimBus53[6]  = s_logisimNet6;
   assign s_logisimBus53[7]  = s_logisimNet3;
   assign s_logisimBus53[8]  = s_logisimNet17;
   assign s_logisimBus53[9]  = s_logisimNet14;
   assign s_logisimBus54[0]  = s_logisimNet40;
   assign s_logisimBus54[10] = s_logisimNet28;
   assign s_logisimBus54[11] = s_logisimNet5;
   assign s_logisimBus54[12] = s_logisimNet32;
   assign s_logisimBus54[13] = s_logisimNet13;
   assign s_logisimBus54[14] = s_logisimNet27;
   assign s_logisimBus54[15] = s_logisimNet6;
   assign s_logisimBus54[16] = s_logisimNet3;
   assign s_logisimBus54[17] = s_logisimNet17;
   assign s_logisimBus54[18] = s_logisimNet14;
   assign s_logisimBus54[19] = s_logisimNet24;
   assign s_logisimBus54[1]  = s_logisimNet46;
   assign s_logisimBus54[20] = s_logisimNet4;
   assign s_logisimBus54[21] = s_logisimNet22;
   assign s_logisimBus54[22] = s_logisimNet21;
   assign s_logisimBus54[23] = s_logisimNet20;
   assign s_logisimBus54[24] = s_logisimNet7;
   assign s_logisimBus54[25] = s_logisimNet2;
   assign s_logisimBus54[26] = s_logisimNet23;
   assign s_logisimBus54[27] = s_logisimNet0;
   assign s_logisimBus54[28] = s_logisimNet19;
   assign s_logisimBus54[29] = s_logisimNet16;
   assign s_logisimBus54[2]  = s_logisimNet37;
   assign s_logisimBus54[30] = s_logisimNet8;
   assign s_logisimBus54[31] = s_logisimNet1;
   assign s_logisimBus54[3]  = s_logisimNet35;
   assign s_logisimBus54[4]  = s_logisimNet44;
   assign s_logisimBus54[5]  = s_logisimNet29;
   assign s_logisimBus54[6]  = s_logisimNet15;
   assign s_logisimBus54[7]  = s_logisimNet34;
   assign s_logisimBus54[8]  = s_logisimNet12;
   assign s_logisimBus54[9]  = s_logisimNet10;
   assign s_logisimBus55[0]  = s_logisimNet12;
   assign s_logisimBus55[10] = s_logisimNet14;
   assign s_logisimBus55[11] = s_logisimNet24;
   assign s_logisimBus55[12] = s_logisimNet4;
   assign s_logisimBus55[13] = s_logisimNet22;
   assign s_logisimBus55[14] = s_logisimNet21;
   assign s_logisimBus55[15] = s_logisimNet20;
   assign s_logisimBus55[16] = s_logisimNet7;
   assign s_logisimBus55[17] = s_logisimNet2;
   assign s_logisimBus55[18] = s_logisimNet23;
   assign s_logisimBus55[19] = s_logisimNet0;
   assign s_logisimBus55[1]  = s_logisimNet10;
   assign s_logisimBus55[20] = s_logisimNet19;
   assign s_logisimBus55[21] = s_logisimNet16;
   assign s_logisimBus55[22] = s_logisimNet8;
   assign s_logisimBus55[23] = s_logisimNet1;
   assign s_logisimBus55[24] = s_logisimNet1;
   assign s_logisimBus55[25] = s_logisimNet1;
   assign s_logisimBus55[26] = s_logisimNet1;
   assign s_logisimBus55[27] = s_logisimNet1;
   assign s_logisimBus55[28] = s_logisimNet1;
   assign s_logisimBus55[29] = s_logisimNet1;
   assign s_logisimBus55[2]  = s_logisimNet28;
   assign s_logisimBus55[30] = s_logisimNet1;
   assign s_logisimBus55[31] = s_logisimNet1;
   assign s_logisimBus55[3]  = s_logisimNet5;
   assign s_logisimBus55[4]  = s_logisimNet32;
   assign s_logisimBus55[5]  = s_logisimNet13;
   assign s_logisimBus55[6]  = s_logisimNet27;
   assign s_logisimBus55[7]  = s_logisimNet6;
   assign s_logisimBus55[8]  = s_logisimNet3;
   assign s_logisimBus55[9]  = s_logisimNet17;
   assign s_logisimBus56[0]  = s_logisimNet17;
   assign s_logisimBus56[10] = s_logisimNet0;
   assign s_logisimBus56[11] = s_logisimNet19;
   assign s_logisimBus56[12] = s_logisimNet16;
   assign s_logisimBus56[13] = s_logisimNet8;
   assign s_logisimBus56[14] = s_logisimNet1;
   assign s_logisimBus56[15] = s_logisimNet1;
   assign s_logisimBus56[16] = s_logisimNet1;
   assign s_logisimBus56[17] = s_logisimNet1;
   assign s_logisimBus56[18] = s_logisimNet1;
   assign s_logisimBus56[19] = s_logisimNet1;
   assign s_logisimBus56[1]  = s_logisimNet14;
   assign s_logisimBus56[20] = s_logisimNet1;
   assign s_logisimBus56[21] = s_logisimNet1;
   assign s_logisimBus56[22] = s_logisimNet1;
   assign s_logisimBus56[23] = s_logisimNet1;
   assign s_logisimBus56[24] = s_logisimNet1;
   assign s_logisimBus56[25] = s_logisimNet1;
   assign s_logisimBus56[26] = s_logisimNet1;
   assign s_logisimBus56[27] = s_logisimNet1;
   assign s_logisimBus56[28] = s_logisimNet1;
   assign s_logisimBus56[29] = s_logisimNet1;
   assign s_logisimBus56[2]  = s_logisimNet24;
   assign s_logisimBus56[30] = s_logisimNet1;
   assign s_logisimBus56[31] = s_logisimNet1;
   assign s_logisimBus56[3]  = s_logisimNet4;
   assign s_logisimBus56[4]  = s_logisimNet22;
   assign s_logisimBus56[5]  = s_logisimNet21;
   assign s_logisimBus56[6]  = s_logisimNet20;
   assign s_logisimBus56[7]  = s_logisimNet7;
   assign s_logisimBus56[8]  = s_logisimNet2;
   assign s_logisimBus56[9]  = s_logisimNet23;
   assign s_logisimBus57[0]  = s_logisimNet20;
   assign s_logisimBus57[10] = s_logisimNet1;
   assign s_logisimBus57[11] = s_logisimNet1;
   assign s_logisimBus57[12] = s_logisimNet1;
   assign s_logisimBus57[13] = s_logisimNet1;
   assign s_logisimBus57[14] = s_logisimNet1;
   assign s_logisimBus57[15] = s_logisimNet1;
   assign s_logisimBus57[16] = s_logisimNet1;
   assign s_logisimBus57[17] = s_logisimNet1;
   assign s_logisimBus57[18] = s_logisimNet1;
   assign s_logisimBus57[19] = s_logisimNet1;
   assign s_logisimBus57[1]  = s_logisimNet7;
   assign s_logisimBus57[20] = s_logisimNet1;
   assign s_logisimBus57[21] = s_logisimNet1;
   assign s_logisimBus57[22] = s_logisimNet1;
   assign s_logisimBus57[23] = s_logisimNet1;
   assign s_logisimBus57[24] = s_logisimNet1;
   assign s_logisimBus57[25] = s_logisimNet1;
   assign s_logisimBus57[26] = s_logisimNet1;
   assign s_logisimBus57[27] = s_logisimNet1;
   assign s_logisimBus57[28] = s_logisimNet1;
   assign s_logisimBus57[29] = s_logisimNet1;
   assign s_logisimBus57[2]  = s_logisimNet2;
   assign s_logisimBus57[30] = s_logisimNet1;
   assign s_logisimBus57[31] = s_logisimNet1;
   assign s_logisimBus57[3]  = s_logisimNet23;
   assign s_logisimBus57[4]  = s_logisimNet0;
   assign s_logisimBus57[5]  = s_logisimNet19;
   assign s_logisimBus57[6]  = s_logisimNet16;
   assign s_logisimBus57[7]  = s_logisimNet8;
   assign s_logisimBus57[8]  = s_logisimNet1;
   assign s_logisimBus57[9]  = s_logisimNet1;
   assign s_logisimBus58[0]  = s_logisimNet44;
   assign s_logisimBus58[10] = s_logisimNet27;
   assign s_logisimBus58[11] = s_logisimNet6;
   assign s_logisimBus58[12] = s_logisimNet3;
   assign s_logisimBus58[13] = s_logisimNet17;
   assign s_logisimBus58[14] = s_logisimNet14;
   assign s_logisimBus58[15] = s_logisimNet24;
   assign s_logisimBus58[16] = s_logisimNet4;
   assign s_logisimBus58[17] = s_logisimNet22;
   assign s_logisimBus58[18] = s_logisimNet21;
   assign s_logisimBus58[19] = s_logisimNet20;
   assign s_logisimBus58[1]  = s_logisimNet29;
   assign s_logisimBus58[20] = s_logisimNet7;
   assign s_logisimBus58[21] = s_logisimNet2;
   assign s_logisimBus58[22] = s_logisimNet23;
   assign s_logisimBus58[23] = s_logisimNet0;
   assign s_logisimBus58[24] = s_logisimNet19;
   assign s_logisimBus58[25] = s_logisimNet16;
   assign s_logisimBus58[26] = s_logisimNet8;
   assign s_logisimBus58[27] = s_logisimNet1;
   assign s_logisimBus58[28] = s_logisimNet1;
   assign s_logisimBus58[29] = s_logisimNet1;
   assign s_logisimBus58[2]  = s_logisimNet15;
   assign s_logisimBus58[30] = s_logisimNet1;
   assign s_logisimBus58[31] = s_logisimNet1;
   assign s_logisimBus58[3]  = s_logisimNet34;
   assign s_logisimBus58[4]  = s_logisimNet12;
   assign s_logisimBus58[5]  = s_logisimNet10;
   assign s_logisimBus58[6]  = s_logisimNet28;
   assign s_logisimBus58[7]  = s_logisimNet5;
   assign s_logisimBus58[8]  = s_logisimNet32;
   assign s_logisimBus58[9]  = s_logisimNet13;
   assign s_logisimBus59[0]  = s_logisimNet3;
   assign s_logisimBus59[10] = s_logisimNet23;
   assign s_logisimBus59[11] = s_logisimNet0;
   assign s_logisimBus59[12] = s_logisimNet19;
   assign s_logisimBus59[13] = s_logisimNet16;
   assign s_logisimBus59[14] = s_logisimNet8;
   assign s_logisimBus59[15] = s_logisimNet1;
   assign s_logisimBus59[16] = s_logisimNet1;
   assign s_logisimBus59[17] = s_logisimNet1;
   assign s_logisimBus59[18] = s_logisimNet1;
   assign s_logisimBus59[19] = s_logisimNet1;
   assign s_logisimBus59[1]  = s_logisimNet17;
   assign s_logisimBus59[20] = s_logisimNet1;
   assign s_logisimBus59[21] = s_logisimNet1;
   assign s_logisimBus59[22] = s_logisimNet1;
   assign s_logisimBus59[23] = s_logisimNet1;
   assign s_logisimBus59[24] = s_logisimNet1;
   assign s_logisimBus59[25] = s_logisimNet1;
   assign s_logisimBus59[26] = s_logisimNet1;
   assign s_logisimBus59[27] = s_logisimNet1;
   assign s_logisimBus59[28] = s_logisimNet1;
   assign s_logisimBus59[29] = s_logisimNet1;
   assign s_logisimBus59[2]  = s_logisimNet14;
   assign s_logisimBus59[30] = s_logisimNet1;
   assign s_logisimBus59[31] = s_logisimNet1;
   assign s_logisimBus59[3]  = s_logisimNet24;
   assign s_logisimBus59[4]  = s_logisimNet4;
   assign s_logisimBus59[5]  = s_logisimNet22;
   assign s_logisimBus59[6]  = s_logisimNet21;
   assign s_logisimBus59[7]  = s_logisimNet20;
   assign s_logisimBus59[8]  = s_logisimNet7;
   assign s_logisimBus59[9]  = s_logisimNet2;
   assign s_logisimBus60[0]  = s_logisimNet22;
   assign s_logisimBus60[10] = s_logisimNet1;
   assign s_logisimBus60[11] = s_logisimNet1;
   assign s_logisimBus60[12] = s_logisimNet1;
   assign s_logisimBus60[13] = s_logisimNet1;
   assign s_logisimBus60[14] = s_logisimNet1;
   assign s_logisimBus60[15] = s_logisimNet1;
   assign s_logisimBus60[16] = s_logisimNet1;
   assign s_logisimBus60[17] = s_logisimNet1;
   assign s_logisimBus60[18] = s_logisimNet1;
   assign s_logisimBus60[19] = s_logisimNet1;
   assign s_logisimBus60[1]  = s_logisimNet21;
   assign s_logisimBus60[20] = s_logisimNet1;
   assign s_logisimBus60[21] = s_logisimNet1;
   assign s_logisimBus60[22] = s_logisimNet1;
   assign s_logisimBus60[23] = s_logisimNet1;
   assign s_logisimBus60[24] = s_logisimNet1;
   assign s_logisimBus60[25] = s_logisimNet1;
   assign s_logisimBus60[26] = s_logisimNet1;
   assign s_logisimBus60[27] = s_logisimNet1;
   assign s_logisimBus60[28] = s_logisimNet1;
   assign s_logisimBus60[29] = s_logisimNet1;
   assign s_logisimBus60[2]  = s_logisimNet20;
   assign s_logisimBus60[30] = s_logisimNet1;
   assign s_logisimBus60[31] = s_logisimNet1;
   assign s_logisimBus60[3]  = s_logisimNet7;
   assign s_logisimBus60[4]  = s_logisimNet2;
   assign s_logisimBus60[5]  = s_logisimNet23;
   assign s_logisimBus60[6]  = s_logisimNet0;
   assign s_logisimBus60[7]  = s_logisimNet19;
   assign s_logisimBus60[8]  = s_logisimNet16;
   assign s_logisimBus60[9]  = s_logisimNet8;
   assign s_logisimBus62[0]  = s_logisimNet7;
   assign s_logisimBus62[10] = s_logisimNet1;
   assign s_logisimBus62[11] = s_logisimNet1;
   assign s_logisimBus62[12] = s_logisimNet1;
   assign s_logisimBus62[13] = s_logisimNet1;
   assign s_logisimBus62[14] = s_logisimNet1;
   assign s_logisimBus62[15] = s_logisimNet1;
   assign s_logisimBus62[16] = s_logisimNet1;
   assign s_logisimBus62[17] = s_logisimNet1;
   assign s_logisimBus62[18] = s_logisimNet1;
   assign s_logisimBus62[19] = s_logisimNet1;
   assign s_logisimBus62[1]  = s_logisimNet2;
   assign s_logisimBus62[20] = s_logisimNet1;
   assign s_logisimBus62[21] = s_logisimNet1;
   assign s_logisimBus62[22] = s_logisimNet1;
   assign s_logisimBus62[23] = s_logisimNet1;
   assign s_logisimBus62[24] = s_logisimNet1;
   assign s_logisimBus62[25] = s_logisimNet1;
   assign s_logisimBus62[26] = s_logisimNet1;
   assign s_logisimBus62[27] = s_logisimNet1;
   assign s_logisimBus62[28] = s_logisimNet1;
   assign s_logisimBus62[29] = s_logisimNet1;
   assign s_logisimBus62[2]  = s_logisimNet23;
   assign s_logisimBus62[30] = s_logisimNet1;
   assign s_logisimBus62[31] = s_logisimNet1;
   assign s_logisimBus62[3]  = s_logisimNet0;
   assign s_logisimBus62[4]  = s_logisimNet19;
   assign s_logisimBus62[5]  = s_logisimNet16;
   assign s_logisimBus62[6]  = s_logisimNet8;
   assign s_logisimBus62[7]  = s_logisimNet1;
   assign s_logisimBus62[8]  = s_logisimNet1;
   assign s_logisimBus62[9]  = s_logisimNet1;
   assign s_logisimBus63[0]  = s_logisimNet35;
   assign s_logisimBus63[10] = s_logisimNet13;
   assign s_logisimBus63[11] = s_logisimNet27;
   assign s_logisimBus63[12] = s_logisimNet6;
   assign s_logisimBus63[13] = s_logisimNet3;
   assign s_logisimBus63[14] = s_logisimNet17;
   assign s_logisimBus63[15] = s_logisimNet14;
   assign s_logisimBus63[16] = s_logisimNet24;
   assign s_logisimBus63[17] = s_logisimNet4;
   assign s_logisimBus63[18] = s_logisimNet22;
   assign s_logisimBus63[19] = s_logisimNet21;
   assign s_logisimBus63[1]  = s_logisimNet44;
   assign s_logisimBus63[20] = s_logisimNet20;
   assign s_logisimBus63[21] = s_logisimNet7;
   assign s_logisimBus63[22] = s_logisimNet2;
   assign s_logisimBus63[23] = s_logisimNet23;
   assign s_logisimBus63[24] = s_logisimNet0;
   assign s_logisimBus63[25] = s_logisimNet19;
   assign s_logisimBus63[26] = s_logisimNet16;
   assign s_logisimBus63[27] = s_logisimNet8;
   assign s_logisimBus63[28] = s_logisimNet1;
   assign s_logisimBus63[29] = s_logisimNet1;
   assign s_logisimBus63[2]  = s_logisimNet29;
   assign s_logisimBus63[30] = s_logisimNet1;
   assign s_logisimBus63[31] = s_logisimNet1;
   assign s_logisimBus63[3]  = s_logisimNet15;
   assign s_logisimBus63[4]  = s_logisimNet34;
   assign s_logisimBus63[5]  = s_logisimNet12;
   assign s_logisimBus63[6]  = s_logisimNet10;
   assign s_logisimBus63[7]  = s_logisimNet28;
   assign s_logisimBus63[8]  = s_logisimNet5;
   assign s_logisimBus63[9]  = s_logisimNet32;
   assign s_logisimBus64[0]  = s_logisimNet4;
   assign s_logisimBus64[10] = s_logisimNet8;
   assign s_logisimBus64[11] = s_logisimNet1;
   assign s_logisimBus64[12] = s_logisimNet1;
   assign s_logisimBus64[13] = s_logisimNet1;
   assign s_logisimBus64[14] = s_logisimNet1;
   assign s_logisimBus64[15] = s_logisimNet1;
   assign s_logisimBus64[16] = s_logisimNet1;
   assign s_logisimBus64[17] = s_logisimNet1;
   assign s_logisimBus64[18] = s_logisimNet1;
   assign s_logisimBus64[19] = s_logisimNet1;
   assign s_logisimBus64[1]  = s_logisimNet22;
   assign s_logisimBus64[20] = s_logisimNet1;
   assign s_logisimBus64[21] = s_logisimNet1;
   assign s_logisimBus64[22] = s_logisimNet1;
   assign s_logisimBus64[23] = s_logisimNet1;
   assign s_logisimBus64[24] = s_logisimNet1;
   assign s_logisimBus64[25] = s_logisimNet1;
   assign s_logisimBus64[26] = s_logisimNet1;
   assign s_logisimBus64[27] = s_logisimNet1;
   assign s_logisimBus64[28] = s_logisimNet1;
   assign s_logisimBus64[29] = s_logisimNet1;
   assign s_logisimBus64[2]  = s_logisimNet21;
   assign s_logisimBus64[30] = s_logisimNet1;
   assign s_logisimBus64[31] = s_logisimNet1;
   assign s_logisimBus64[3]  = s_logisimNet20;
   assign s_logisimBus64[4]  = s_logisimNet7;
   assign s_logisimBus64[5]  = s_logisimNet2;
   assign s_logisimBus64[6]  = s_logisimNet23;
   assign s_logisimBus64[7]  = s_logisimNet0;
   assign s_logisimBus64[8]  = s_logisimNet19;
   assign s_logisimBus64[9]  = s_logisimNet16;
   assign s_logisimBus65[0]  = s_logisimNet27;
   assign s_logisimBus65[10] = s_logisimNet7;
   assign s_logisimBus65[11] = s_logisimNet2;
   assign s_logisimBus65[12] = s_logisimNet23;
   assign s_logisimBus65[13] = s_logisimNet0;
   assign s_logisimBus65[14] = s_logisimNet19;
   assign s_logisimBus65[15] = s_logisimNet16;
   assign s_logisimBus65[16] = s_logisimNet8;
   assign s_logisimBus65[17] = s_logisimNet1;
   assign s_logisimBus65[18] = s_logisimNet1;
   assign s_logisimBus65[19] = s_logisimNet1;
   assign s_logisimBus65[1]  = s_logisimNet6;
   assign s_logisimBus65[20] = s_logisimNet1;
   assign s_logisimBus65[21] = s_logisimNet1;
   assign s_logisimBus65[22] = s_logisimNet1;
   assign s_logisimBus65[23] = s_logisimNet1;
   assign s_logisimBus65[24] = s_logisimNet1;
   assign s_logisimBus65[25] = s_logisimNet1;
   assign s_logisimBus65[26] = s_logisimNet1;
   assign s_logisimBus65[27] = s_logisimNet1;
   assign s_logisimBus65[28] = s_logisimNet1;
   assign s_logisimBus65[29] = s_logisimNet1;
   assign s_logisimBus65[2]  = s_logisimNet3;
   assign s_logisimBus65[30] = s_logisimNet1;
   assign s_logisimBus65[31] = s_logisimNet1;
   assign s_logisimBus65[3]  = s_logisimNet17;
   assign s_logisimBus65[4]  = s_logisimNet14;
   assign s_logisimBus65[5]  = s_logisimNet24;
   assign s_logisimBus65[6]  = s_logisimNet4;
   assign s_logisimBus65[7]  = s_logisimNet22;
   assign s_logisimBus65[8]  = s_logisimNet21;
   assign s_logisimBus65[9]  = s_logisimNet20;
   assign s_logisimNet0      = s_logisimBus25[28];
   assign s_logisimNet10     = s_logisimBus25[10];
   assign s_logisimNet12     = s_logisimBus25[9];
   assign s_logisimNet13     = s_logisimBus25[14];
   assign s_logisimNet14     = s_logisimBus25[19];
   assign s_logisimNet15     = s_logisimBus25[7];
   assign s_logisimNet16     = s_logisimBus25[30];
   assign s_logisimNet17     = s_logisimBus25[18];
   assign s_logisimNet19     = s_logisimBus25[29];
   assign s_logisimNet2      = s_logisimBus25[26];
   assign s_logisimNet20     = s_logisimBus25[24];
   assign s_logisimNet21     = s_logisimBus25[23];
   assign s_logisimNet22     = s_logisimBus25[22];
   assign s_logisimNet23     = s_logisimBus25[27];
   assign s_logisimNet24     = s_logisimBus25[20];
   assign s_logisimNet27     = s_logisimBus25[15];
   assign s_logisimNet28     = s_logisimBus25[11];
   assign s_logisimNet29     = s_logisimBus25[6];
   assign s_logisimNet3      = s_logisimBus25[17];
   assign s_logisimNet32     = s_logisimBus25[13];
   assign s_logisimNet34     = s_logisimBus25[8];
   assign s_logisimNet35     = s_logisimBus25[4];
   assign s_logisimNet37     = s_logisimBus25[3];
   assign s_logisimNet4      = s_logisimBus25[21];
   assign s_logisimNet40     = s_logisimBus25[1];
   assign s_logisimNet44     = s_logisimBus25[5];
   assign s_logisimNet46     = s_logisimBus25[2];
   assign s_logisimNet5      = s_logisimBus25[12];
   assign s_logisimNet6      = s_logisimBus25[16];
   assign s_logisimNet7      = s_logisimBus25[25];
   assign s_logisimNet8      = s_logisimBus25[31];

   /*******************************************************************************
   ** Here all input connections are defined                                     **
   *******************************************************************************/
   assign s_logisimBus25[31:0] = in1;
   assign s_logisimBus9[4:0]   = shift;

   /*******************************************************************************
   ** Here all output connections are defined                                    **
   *******************************************************************************/
   assign out1 = s_logisimBus61[31:0];

   /*******************************************************************************
   ** Here all in-lined components are defined                                   **
   *******************************************************************************/

   // Constant
   assign  s_logisimNet1  =  1'b0;


   /*******************************************************************************
   ** Here all normal components are defined                                     **
   *******************************************************************************/
   Multiplexer_bus_32 #(.nrOfBits(32))
      PLEXERS_1 (.enable(1'b1),
                 .muxIn_0(s_logisimBus25[31:0]),
                 .muxIn_1(s_logisimBus54[31:0]),
                 .muxIn_10(s_logisimBus53[31:0]),
                 .muxIn_11(s_logisimBus39[31:0]),
                 .muxIn_12(s_logisimBus33[31:0]),
                 .muxIn_13(s_logisimBus18[31:0]),
                 .muxIn_14(s_logisimBus47[31:0]),
                 .muxIn_15(s_logisimBus65[31:0]),
                 .muxIn_16(s_logisimBus52[31:0]),
                 .muxIn_17(s_logisimBus59[31:0]),
                 .muxIn_18(s_logisimBus56[31:0]),
                 .muxIn_19(s_logisimBus42[31:0]),
                 .muxIn_2(s_logisimBus11[31:0]),
                 .muxIn_20(s_logisimBus36[31:0]),
                 .muxIn_21(s_logisimBus64[31:0]),
                 .muxIn_22(s_logisimBus60[31:0]),
                 .muxIn_23(s_logisimBus50[31:0]),
                 .muxIn_24(s_logisimBus57[31:0]),
                 .muxIn_25(s_logisimBus62[31:0]),
                 .muxIn_26(s_logisimBus43[31:0]),
                 .muxIn_27(s_logisimBus49[31:0]),
                 .muxIn_28(s_logisimBus30[31:0]),
                 .muxIn_29(s_logisimBus31[31:0]),
                 .muxIn_3(s_logisimBus26[31:0]),
                 .muxIn_30(s_logisimBus38[31:0]),
                 .muxIn_31(s_logisimBus48[31:0]),
                 .muxIn_4(s_logisimBus63[31:0]),
                 .muxIn_5(s_logisimBus58[31:0]),
                 .muxIn_6(s_logisimBus45[31:0]),
                 .muxIn_7(s_logisimBus41[31:0]),
                 .muxIn_8(s_logisimBus51[31:0]),
                 .muxIn_9(s_logisimBus55[31:0]),
                 .muxOut(s_logisimBus61[31:0]),
                 .sel(s_logisimBus9[4:0]));


endmodule
